library verilog;
use verilog.vl_types.all;
entity BT3_vlg_vec_tst is
end BT3_vlg_vec_tst;
