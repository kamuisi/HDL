library verilog;
use verilog.vl_types.all;
entity moore_vlg_vec_tst is
end moore_vlg_vec_tst;
