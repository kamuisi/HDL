module full_adder_4bit_0(A, B, Cin, S, Cout);
input [3:0] A, B;
input Cin;
output [3:0] S;
output Cout;
wire w0, w1, w2;

full_adder (A[0], B[0], Cin, S[0], w0);
full_adder (A[1], B[1], w0, S[1], w1);
full_adder (A[2], A[2], w1, S[2], w2);
full_adder (A[3], A[3], w2, S[3], Cout);

endmodule