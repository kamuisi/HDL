library verilog;
use verilog.vl_types.all;
entity lifo_stack_tb is
end lifo_stack_tb;
