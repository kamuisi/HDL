library verilog;
use verilog.vl_types.all;
entity CLA_3b_vlg_vec_tst is
end CLA_3b_vlg_vec_tst;
