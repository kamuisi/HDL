module full_adder_4bit_2(A, B, Cin, S, Cout);
input [3:0] A, B;
input Cin;
output reg [3:0] S;
output reg Cout;

always @(*)
	begin
		{Cout, S} <= A + B + Cin;
	end
endmodule	