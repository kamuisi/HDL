library verilog;
use verilog.vl_types.all;
entity full_adder_4bit_0_vlg_check_tst is
    port(
        Cout            : in     vl_logic;
        S               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end full_adder_4bit_0_vlg_check_tst;
