library verilog;
use verilog.vl_types.all;
entity mealy_vlg_vec_tst is
end mealy_vlg_vec_tst;
