library verilog;
use verilog.vl_types.all;
entity SRAM_vlg_vec_tst is
end SRAM_vlg_vec_tst;
