library verilog;
use verilog.vl_types.all;
entity lab_2_1_vlg_vec_tst is
end lab_2_1_vlg_vec_tst;
