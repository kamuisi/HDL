library verilog;
use verilog.vl_types.all;
entity BT6_tb is
end BT6_tb;
